-------------------------------------------
-- Block code:  dds_top.vhd
-- History: 	20.Apr.2018 - 1st version (Felipe Tanios)
--                 
-- Function: Top for direct digital synthesis block
------------------------------------------- 

-- Library & Use Statements
LIBRARY ieee;
use ieee.std_logic_1164.all;
LIBRARY work;
USE work.tone_gen_pkg.all;

entity dds_top is
	port(
		tone_cmd		: in    std_logic_vector(1 downto 0);
		wave_ctrl		: in 	std_logic_vector(1 downto 0);
		clock			: in    std_logic;
		strobe_i		: in 	  std_logic;
		rst_n			: in    std_logic;
		dacdat_g_out	: out 	std_logic_vector(N_AUDIO - 1 downto 0)
	);
end dds_top;

ARCHITECTURE struct OF dds_top IS

	SIGNAL top_phi_incr 	: std_logic_vector(N_CUM-1 downto 0);
	SIGNAL top_tone_on  	: std_logic;

	COMPONENT tone_decoder is
        port(
			tone_cmd_i		: in	std_logic_vector(1 downto 0);
			phi_incr_o		: out 	std_logic_vector(N_CUM-1 downto 0);
			tone_on_o		: out	std_logic
        );
	end COMPONENT;
	
	COMPONENT DDS is
		port(
			tone_on_i		: in    std_logic;
			phi_incr_i		: in    std_logic_vector(N_CUM-1 downto 0);
			strobe_in		: in    std_logic;
			clk, reset_n	: in	std_logic;
			wave_i			: in 	std_logic_vector(1 downto 0);
			dacdat_g_o		: out 	std_logic_vector(N_AUDIO - 1 downto 0)
		);
	end COMPONENT;
	
	BEGIN
	
		inst_tone_decoder: tone_decoder
        port map(
			tone_cmd_i		=> tone_cmd,
			phi_incr_o		=> top_phi_incr,
			tone_on_o		=> top_tone_on
        );
	
		inst_dds: DDS
		port map(
			tone_on_i		=> top_tone_on,
			phi_incr_i		=> top_phi_incr,
			strobe_in		=> strobe_i,
			clk				=> clock,
			reset_n			=> rst_n,
			wave_i			=> wave_ctrl,
			dacdat_g_o		=> dacdat_g_out
		);

END struct;	